-------------------------------------------------------------------------------
-- Title      : COMP.CE.240, Exercise 12
-- Project    : 
-------------------------------------------------------------------------------
-- File       : tb_i2c_config.vhd
-- Author     : Group 21, Kaakkolammi Henrik, xxx xxx
-- Company    : 
-- Created    : 2021-02-21
-- Last update: 2021-02-21
-- Platform   : 
-- Standard   : VHDL'93/02
-------------------------------------------------------------------------------
-- Description: I2C controller testbench
-------------------------------------------------------------------------------
-- Copyright (c) 2021
-------------------------------------------------------------------------------
-- Revisions  :
-- Date        Version  Author      Description
-- 2021-02-21  1.0      Kaakkolammi Created
-------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;

-------------------------------------------------------------------------------
-- Empty entity
-------------------------------------------------------------------------------

entity tb_i2c_config is
end tb_i2c_config;

-------------------------------------------------------------------------------
-- Architecture
-------------------------------------------------------------------------------
architecture testbench of tb_i2c_config is

  -- Number of parameters to expect
  constant n_params_c     : integer := 15;
  constant n_leds_c       : integer := 4;
  constant i2c_freq_c     : integer := 20000;
  constant ref_freq_c     : integer := 50000000;
  constant clock_period_c : time    := 20 ns;

  -- Every transmission consists several bytes and every byte contains given
  -- amount of bits. 
  constant n_bytes_c       : integer := 3;
  constant bit_count_max_c : integer := 8;

  -- Signals fed to the DUV
  signal clk   : std_logic := '0';  -- Remember that default values supported
  signal rst_n : std_logic := '0';      -- only in synthesis

  -- The DUV prototype
  component i2c_config
    generic (
      ref_clk_freq_g : integer;
      i2c_freq_g     : integer;
      n_params_g     : integer;
	    n_leds_g       : integer);
    port (
      clk              : in    std_logic;
      rst_n            : in    std_logic;
      sdat_inout       : inout std_logic;
      sclk_out         : out   std_logic;
      param_status_out : out   std_logic_vector(n_leds_g-1 downto 0);
      finished_out     : out   std_logic
      );
  end component;

  -- Signals coming from the DUV
  signal sdat         : std_logic := 'Z';
  signal sclk         : std_logic;
  signal param_status : std_logic_vector(n_leds_c-1 downto 0);
  signal finished     : std_logic;

  -- To hold the value that will be driven to sdat when sclk is high.
  signal sdat_r : std_logic;

  -- Counters for receiving bits and bytes
  signal bit_counter_r  : integer range 0 to bit_count_max_c-1;
  signal byte_counter_r : integer range 0 to n_bytes_c-1;

  -- States for the FSM
  type   states is (wait_start, read_byte, send_ack, wait_stop);
  signal curr_state_r : states;

  -- Previous values of the I2C signals for edge detection
  signal sdat_old_r : std_logic;
  signal sclk_old_r : std_logic;

  -- Data storages for transfers
  signal sdat_byte_r          : std_logic_vector(bit_count_max_c-1 downto 0);
  signal sdat_transfer_r      : std_logic_vector(
                                bit_count_max_c*n_bytes_c-1 downto 0);
  signal sdat_byte_counter_r  : integer range 0 to n_bytes_c-1;
  
  -- Flag for NACK
  signal sdat_nack_r        : std_logic;
  signal sdat_nack_tested_r : std_logic;

  -- All the other data to send is in the following array:
  type data_array is array (n_params_c-1 downto 0) of std_logic_vector(15 DOWNTO 0);
  signal i2c_data_array_r : data_array;
  -- Flag array to keep track of which commands have been received
  signal i2c_data_flags_r : std_logic_vector(n_params_c-1 downto 0);
  -- Flag for unrecognised configuration data received
  signal unknown_config_data_r : std_logic;

begin  -- testbench

  i2c_data_array_r(0) <= "0001110110000000";
  i2c_data_array_r(1) <= "0010011100000100";
  i2c_data_array_r(2) <= "0010001000001011";
  i2c_data_array_r(3) <= "0010100000000000";
  i2c_data_array_r(4) <= "0010100110000001";
  i2c_data_array_r(5) <= "0110100100001000";
  i2c_data_array_r(6) <= "0110101000000000";
  i2c_data_array_r(7) <= "0100011111100001";
  i2c_data_array_r(8) <= "0110101100001001";
  i2c_data_array_r(9) <= "0110110000001000";
  i2c_data_array_r(10) <= "0100101100001000";
  i2c_data_array_r(11) <= "0100110000001000";
  i2c_data_array_r(12) <= "0110111010001000";
  i2c_data_array_r(13) <= "0110111110001000";
  i2c_data_array_r(14) <= "0101000111110001";

  clk   <= not clk after clock_period_c/2;
  rst_n <= '1'     after clock_period_c*4;

  -- Assign sdat_r when sclk is active, otherwise 'Z'.
  -- Note that sdat_r is usually 'Z'
  with sclk select
    sdat <=
        sdat_r when '1',
        'Z'    when others;


  -- Component instantiation
  i2c_config_1 : i2c_config
    generic map (
      ref_clk_freq_g => ref_freq_c,
      i2c_freq_g     => i2c_freq_c,
      n_params_g     => n_params_c,
	    n_leds_g => n_leds_c)
    port map (
      clk              => clk,
      rst_n            => rst_n,
      sdat_inout       => sdat,
      sclk_out         => sclk,
      param_status_out => param_status,
      finished_out     => finished);

  -----------------------------------------------------------------------------
  -- The main process that controls the behavior of the test bench
  fsm_proc : process (clk, rst_n)
  begin  -- process fsm_proc
    if rst_n = '0' then                 -- asynchronous reset (active low)

      curr_state_r <= wait_start;

      sdat_old_r <= '0';
      sclk_old_r <= '0';

      byte_counter_r <= 0;
      bit_counter_r  <= 0;

      sdat_r <= 'Z';

      sdat_byte_r <= (others => '0');
      sdat_transfer_r <= (others => '0');
      sdat_byte_counter_r <= 0;

      sdat_nack_r <= '0';
      sdat_nack_tested_r <= '0';

      i2c_data_flags_r <= (others => '0');
      unknown_config_data_r <= '0';
      
    elsif clk'event and clk = '1' then  -- rising clock edge
      -- The previous values are required for the edge detection
      sclk_old_r <= sclk;
      sdat_old_r <= sdat;

      -- Falling edge detection for acknowledge control
      -- Must be done on the falling edge in order to be stable during
      -- the high period of sclk
      if sclk = '0' and sclk_old_r = '1' then
        -- If we are supposed to send ack
        if curr_state_r = send_ack then
          -- Send ack (low = ACK, high = NACK)
          if sdat_nack_r = '0' then
            sdat_r <= '0';
          else
            sdat_r <= '1';
            -- Reset nack back to 0 after testing it
            sdat_nack_r <= '0';
          end if;
        else
          -- Otherwise, sdat is in high impedance state.
          sdat_r <= 'Z';
        end if;
        
      end if;


      -------------------------------------------------------------------------
      -- FSM
      case curr_state_r is
        -----------------------------------------------------------------------
        -- Wait for the start condition
        when wait_start =>
          -- While clk stays high, the sdat falls
          if sclk = '1' and sclk_old_r = '1' and
            sdat_old_r = '1' and sdat = '0' then

            curr_state_r <= read_byte;
          end if;

          --------------------------------------------------------------------
          -- Wait for a byte to be read
        when read_byte =>
          -- Detect a rising edge
          if sclk = '1' and sclk_old_r = '0' then
            -- Save bits
            sdat_byte_r(bit_counter_r) <= sdat;
            -- Indexing down from 23 to 0
            sdat_transfer_r(bit_count_max_c*n_bytes_c-1 - 
              (sdat_byte_counter_r*bit_count_max_c + bit_counter_r)) <= sdat;

            if bit_counter_r /= bit_count_max_c-1 then
              -- Normally just receive a bit
              bit_counter_r <= bit_counter_r + 1;
            else
              -- Byte counter
              if sdat_byte_counter_r = 2 then
                sdat_byte_counter_r <= 0;

                -- Check here if the message is correct
                -- Device address and R/W test
                assert sdat_transfer_r(23 downto 16) = "00110100" report 
                "Incorrect device address" severity failure;

                              
                -- Check configuration values
                -- Asserted at the end of the test
                -- Stays as 1 if no config was found. TODO: Check if assert works
                unknown_config_data_r <= '1';
                for i in 0 to 14 loop
                  if sdat_transfer_r(15 downto 0) = i2c_data_array_r(i) then
                    i2c_data_flags_r(i) <= '1';
                    unknown_config_data_r <= '0';
                  end if;
                end loop;
              else
                sdat_byte_counter_r <= sdat_byte_counter_r + 1;
              end if;

              -- Test NACK by setting sdat_nack_r=1
              -- Will be done once when transfer has arbitrary bit set 1
              if sdat_transfer_r(3) = '1' and sdat_nack_tested_r = '0' then
                sdat_nack_r <= '1';
                sdat_nack_tested_r <= '1';
              end if;

              -- When terminal count is reached, let's send the ack
              curr_state_r  <= send_ack;
              bit_counter_r <= 0;
            end if;  -- Bit counter terminal count
          end if;  -- sclk rising clock edge

          --------------------------------------------------------------------
          -- Send acknowledge
        when send_ack =>
          -- Detect a rising edge
          if sclk = '1' and sclk_old_r = '0' then
            if byte_counter_r /= n_bytes_c-1 then
              -- Transmission continues
              byte_counter_r <= byte_counter_r + 1;
              curr_state_r   <= read_byte;
            else
              -- Transmission is about to stop
              byte_counter_r <= 0;
              curr_state_r   <= wait_stop;
            end if;
          end if;

          ---------------------------------------------------------------------
          -- Wait for the stop condition
        when wait_stop =>
          -- Stop condition detection: sdat rises while sclk stays high
          if sclk = '1' and sclk_old_r = '1' and
            sdat_old_r = '0' and sdat = '1' then

            curr_state_r <= wait_start;
          end if;
      end case;
    end if;
  end process fsm_proc;

  -----------------------------------------------------------------------------
  -- Asserts for verification
  -----------------------------------------------------------------------------

  -- SDAT should never contain X:s.
  assert sdat /= 'X' report "Three state bus in state X" severity failure;
  -- All configurations received should be on the list
  assert rst_n = '0' or unknown_config_data_r = '0' report
    "Unknown configuration received" severity failure;
  
  -- All configs received
  assert rst_n='0' or finished = '0' or i2c_data_flags_r = "111111111111111" report
    "All configurations were not received" severity failure;
  -- End of simulation, but not during the reset
  assert finished = '0' or rst_n = '0' report
    "Simulation done" severity failure;
  
end testbench;
